LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY store_buff IS
	PORT(		
				clock, reset				: IN 	STD_LOGIC; --clock on which to add items
				incoming_indicator		: IN	STD_LOGIC;
				incoming_instruction		: IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
				incoming_address			: IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
				MEM_busy						: IN  STD_LOGIC;
				opcode_out					: OUT STD_LOGIC_VECTOR( 5 DOWNTO 0);
				addr_out						: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
				store_buff_full			: OUT STD_LOGIC := '0';
				store_buff_empty			: OUT STD_LOGIC;
				load_buff_full				: OUT STD_LOGIC := '0';
				ld								: OUT	STD_LOGIC;
				st								: OUT	STD_LOGIC;
				op_code						: OUT STD_LOGIC_VECTOR( 5 DOWNTO 0);
				tester						: OUT STD_LOGIC
		 );
END store_buff;

ARCHITECTURE behavior OF store_buff IS
	
TYPE entry IS
	RECORD
		opcode						: STD_LOGIC_VECTOR( 5 DOWNTO 0); -- 0
		address						: STD_LOGIC_VECTOR(31 DOWNTO 0); -- 1
		isEmpty						: STD_LOGIC;					 		-- 2
	END RECORD;

TYPE store_buff IS ARRAY (0 TO 31) OF entry;

SIGNAL store_buffer	:		store_buff;

TYPE load_buff IS ARRAY (0 TO 31) OF entry;

SIGNAL load_buffer	:		load_buff;

SIGNAL op							:	STD_LOGIC_VECTOR( 5 DOWNTO 0);
SIGNAL addr							:	STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL hold							:  STD_LOGIC;
SIGNAL store_buff_empty_sig	:	STD_LOGIC;
SIGNAL load_in						: 	STD_LOGIC;
SIGNAL store_in					:	STD_LOGIC;

BEGIN
	op 	<= incoming_instruction(31 DOWNTO 26);
	addr	<= incoming_address;
	tester <= store_buffer(31).isEmpty;
	op_code <= op;
	
	ld		<= load_in;
	st		<= store_in;
	
	PROCESS(clock, reset, op, addr, store_buffer, load_buffer, store_buff_empty_sig)
	BEGIN
		IF(reset = '0') THEN
		ELSIF(RISING_EDGE(clock)) THEN
			IF(incoming_indicator = '1') THEN
				IF(op = "100011") THEN -- this is a store
					IF(store_buffer(0).isEmpty = '0') THEN
						store_buffer(0).opcode 	<= op;
						store_buffer(0).address <= addr;
						store_buffer(0).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(1).isEmpty = '0') THEN
						store_buffer(1).opcode 	<= op;
						store_buffer(1).address <= addr;
						store_buffer(1).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(2).isEmpty = '0') THEN
						store_buffer(2).opcode 	<= op;
						store_buffer(2).address <= addr;
						store_buffer(2).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(3).isEmpty = '0') THEN
						store_buffer(3).opcode 	<= op;
						store_buffer(3).address <= addr;
						store_buffer(3).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(4).isEmpty = '0') THEN
						store_buffer(4).opcode 	<= op;
						store_buffer(4).address <= addr;
						store_buffer(4).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(5).isEmpty = '0') THEN
						store_buffer(5).opcode 	<= op;
						store_buffer(5).address <= addr;
						store_buffer(5).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(6).isEmpty = '0') THEN
						store_buffer(6).opcode 	<= op;
						store_buffer(6).address <= addr;
						store_buffer(6).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(7).isEmpty = '0') THEN
						store_buffer(7).opcode 	<= op;
						store_buffer(7).address <= addr;
						store_buffer(7).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(8).isEmpty = '0') THEN
						store_buffer(8).opcode 	<= op;
						store_buffer(8).address <= addr;
						store_buffer(8).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(9).isEmpty = '0') THEN
						store_buffer(9).opcode 	<= op;
						store_buffer(9).address <= addr;
						store_buffer(9).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(10).isEmpty = '0') THEN
						store_buffer(10).opcode 	<= op;
						store_buffer(10).address <= addr;
						store_buffer(10).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(11).isEmpty = '0') THEN
						store_buffer(11).opcode 	<= op;
						store_buffer(11).address <= addr;
						store_buffer(11).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(12).isEmpty = '0') THEN
						store_buffer(12).opcode 	<= op;
						store_buffer(12).address <= addr;
						store_buffer(12).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(13).isEmpty = '0') THEN
						store_buffer(13).opcode 	<= op;
						store_buffer(13).address <= addr;
						store_buffer(13).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(14).isEmpty = '0') THEN
						store_buffer(14).opcode 	<= op;
						store_buffer(14).address <= addr;
						store_buffer(14).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(15).isEmpty = '0') THEN
						store_buffer(15).opcode 	<= op;
						store_buffer(15).address <= addr;
						store_buffer(15).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(16).isEmpty = '0') THEN
						store_buffer(16).opcode 	<= op;
						store_buffer(16).address <= addr;
						store_buffer(16).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(17).isEmpty = '0') THEN
						store_buffer(17).opcode 	<= op;
						store_buffer(17).address <= addr;
						store_buffer(17).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(18).isEmpty = '0') THEN
						store_buffer(18).opcode 	<= op;
						store_buffer(18).address <= addr;
						store_buffer(18).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(19).isEmpty = '0') THEN
						store_buffer(19).opcode 	<= op;
						store_buffer(19).address <= addr;
						store_buffer(19).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(20).isEmpty = '0') THEN
						store_buffer(20).opcode 	<= op;
						store_buffer(20).address <= addr;
						store_buffer(20).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(21).isEmpty = '0') THEN
						store_buffer(21).opcode 	<= op;
						store_buffer(21).address <= addr;
						store_buffer(21).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(22).isEmpty = '0') THEN
						store_buffer(22).opcode 	<= op;
						store_buffer(22).address <= addr;
						store_buffer(22).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(23).isEmpty = '0') THEN
						store_buffer(23).opcode 	<= op;
						store_buffer(23).address <= addr;
						store_buffer(23).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(23).isEmpty = '0') THEN
						store_buffer(23).opcode 	<= op;
						store_buffer(23).address <= addr;
						store_buffer(23).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(24).isEmpty = '0') THEN
						store_buffer(24).opcode 	<= op;
						store_buffer(24).address <= addr;
						store_buffer(24).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(25).isEmpty = '0') THEN
						store_buffer(25).opcode 	<= op;
						store_buffer(25).address <= addr;
						store_buffer(25).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(26).isEmpty = '0') THEN
						store_buffer(26).opcode 	<= op;
						store_buffer(26).address <= addr;
						store_buffer(26).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(27).isEmpty = '0') THEN
						store_buffer(27).opcode 	<= op;
						store_buffer(27).address <= addr;
						store_buffer(27).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(28).isEmpty = '0') THEN
						store_buffer(28).opcode 	<= op;
						store_buffer(28).address <= addr;
						store_buffer(28).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(29).isEmpty = '0') THEN
						store_buffer(29).opcode 	<= op;
						store_buffer(29).address <= addr;
						store_buffer(29).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(30).isEmpty = '0') THEN
						store_buffer(30).opcode 	<= op;
						store_buffer(30).address <= addr;
						store_buffer(30).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSIF(store_buffer(31).isEmpty = '0') THEN
						store_buffer(31).opcode 	<= op;
						store_buffer(31).address <= addr;
						store_buffer(31).isEmpty <= '1';
						--store_buff_full			<= '0';
					ELSE
						--store_buff_full			<= '1';
					END IF;
				ELSIF(op = "101011") THEN -- this is a load
					IF(store_buffer(0).isEmpty = '0') THEN
						load_buffer(0).opcode 	<= op;
						load_buffer(0).address <= addr;
						load_buffer(0).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(1).isEmpty = '0') THEN
						load_buffer(1).opcode 	<= op;
						load_buffer(1).address <= addr;
						load_buffer(1).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(2).isEmpty = '0') THEN
						load_buffer(2).opcode 	<= op;
						load_buffer(2).address <= addr;
						load_buffer(2).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(3).isEmpty = '0') THEN
						load_buffer(3).opcode 	<= op;
						load_buffer(3).address <= addr;
						load_buffer(3).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(4).isEmpty = '0') THEN
						load_buffer(4).opcode 	<= op;
						load_buffer(4).address <= addr;
						load_buffer(4).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(5).isEmpty = '0') THEN
						load_buffer(5).opcode 	<= op;
						load_buffer(5).address <= addr;
						load_buffer(5).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(6).isEmpty = '0') THEN
						load_buffer(6).opcode 	<= op;
						load_buffer(6).address <= addr;
						load_buffer(6).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(7).isEmpty = '0') THEN
						load_buffer(7).opcode 	<= op;
						load_buffer(7).address <= addr;
						load_buffer(7).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(8).isEmpty = '0') THEN
						load_buffer(8).opcode 	<= op;
						load_buffer(8).address <= addr;
						load_buffer(8).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(9).isEmpty = '0') THEN
						load_buffer(9).opcode 	<= op;
						load_buffer(9).address <= addr;
						load_buffer(9).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(10).isEmpty = '0') THEN
						load_buffer(10).opcode 	<= op;
						load_buffer(10).address <= addr;
						load_buffer(10).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(11).isEmpty = '0') THEN
						load_buffer(11).opcode 	<= op;
						load_buffer(11).address <= addr;
						load_buffer(11).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(12).isEmpty = '0') THEN
						load_buffer(12).opcode 	<= op;
						load_buffer(12).address <= addr;
						load_buffer(12).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(13).isEmpty = '0') THEN
						load_buffer(13).opcode 	<= op;
						load_buffer(13).address <= addr;
						load_buffer(13).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(14).isEmpty = '0') THEN
						load_buffer(14).opcode 	<= op;
						load_buffer(14).address <= addr;
						load_buffer(14).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(15).isEmpty = '0') THEN
						load_buffer(15).opcode 	<= op;
						load_buffer(15).address <= addr;
						load_buffer(15).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(16).isEmpty = '0') THEN
						load_buffer(16).opcode 	<= op;
						load_buffer(16).address <= addr;
						load_buffer(16).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(17).isEmpty = '0') THEN
						load_buffer(17).opcode 	<= op;
						load_buffer(17).address <= addr;
						load_buffer(17).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(18).isEmpty = '0') THEN
						load_buffer(18).opcode 	<= op;
						load_buffer(18).address <= addr;
						load_buffer(18).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(19).isEmpty = '0') THEN
						load_buffer(19).opcode 	<= op;
						load_buffer(19).address <= addr;
						load_buffer(19).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(20).isEmpty = '0') THEN
						load_buffer(20).opcode 	<= op;
						load_buffer(20).address <= addr;
						load_buffer(20).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(21).isEmpty = '0') THEN
						load_buffer(21).opcode 	<= op;
						load_buffer(21).address <= addr;
						load_buffer(21).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(22).isEmpty = '0') THEN
						load_buffer(22).opcode 	<= op;
						load_buffer(22).address <= addr;
						load_buffer(22).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(23).isEmpty = '0') THEN
						load_buffer(23).opcode 	<= op;
						load_buffer(23).address <= addr;
						load_buffer(23).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(23).isEmpty = '0') THEN
						load_buffer(23).opcode 	<= op;
						load_buffer(23).address <= addr;
						load_buffer(23).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(24).isEmpty = '0') THEN
						load_buffer(24).opcode 	<= op;
						load_buffer(24).address <= addr;
						load_buffer(24).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(25).isEmpty = '0') THEN
						load_buffer(25).opcode 	<= op;
						load_buffer(25).address <= addr;
						load_buffer(25).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(26).isEmpty = '0') THEN
						load_buffer(26).opcode 	<= op;
						load_buffer(26).address <= addr;
						load_buffer(26).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(27).isEmpty = '0') THEN
						load_buffer(27).opcode 	<= op;
						load_buffer(27).address <= addr;
						load_buffer(27).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(28).isEmpty = '0') THEN
						load_buffer(28).opcode 	<= op;
						load_buffer(28).address <= addr;
						load_buffer(28).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSIF(load_buffer(29).isEmpty = '0') THEN
						load_buffer(29).opcode 	<= op;
						load_buffer(29).address <= addr;
						load_buffer(29).isEmpty <= '1';
						----load_buff_full			<= '0';
					ELSIF(load_buffer(30).isEmpty = '0') THEN
						load_buffer(30).opcode 	<= op;
						load_buffer(30).address <= addr;
						load_buffer(30).isEmpty <= '1';
						----load_buff_full			<= '0';
					ELSIF(load_buffer(31).isEmpty = '0') THEN
						load_buffer(31).opcode 	<= op;
						load_buffer(31).address <= addr;
						load_buffer(31).isEmpty <= '1';
						--load_buff_full			<= '0';
					ELSE
						--load_buff_full			<= '1';
					END IF;
				END IF;
			END IF;
		---
			IF(MEM_busy = '0') THEN--pushing items into the mem unit
				store_in <= '1';
				IF(store_buffer(0).isEmpty = '1') THEN
					addr_out <= store_buffer(0).address;
					opcode_out <= store_buffer(0).opcode;
					store_buffer(0).isEmpty <= '0';
				ELSIF(store_buffer(1).isEmpty = '1') THEN
					addr_out <= store_buffer(1).address;
					opcode_out <= store_buffer(1).opcode;
					store_buffer(1).isEmpty <= '0';
				ELSIF(store_buffer(2).isEmpty = '1') THEN
					addr_out <= store_buffer(2).address;
					opcode_out <= store_buffer(2).opcode;
					store_buffer(2).isEmpty <= '0';
				ELSIF(store_buffer(3).isEmpty = '1') THEN
					addr_out <= store_buffer(3).address;
					opcode_out <= store_buffer(3).opcode;
					store_buffer(3).isEmpty <= '0';
				ELSIF(store_buffer(4).isEmpty = '1') THEN
					addr_out <= store_buffer(4).address;
					opcode_out <= store_buffer(4).opcode;
					store_buffer(4).isEmpty <= '0';
				ELSIF(store_buffer(5).isEmpty = '1') THEN
					addr_out <= store_buffer(5).address;
					opcode_out <= store_buffer(5).opcode;
					store_buffer(5).isEmpty <= '0';
				ELSIF(store_buffer(6).isEmpty = '1') THEN
					addr_out <= store_buffer(6).address;
					opcode_out <= store_buffer(6).opcode;
					store_buffer(6).isEmpty <= '0';
				ELSIF(store_buffer(7).isEmpty = '1') THEN
					addr_out <= store_buffer(7).address;
					opcode_out <= store_buffer(7).opcode;
					store_buffer(7).isEmpty <= '0';
				ELSIF(store_buffer(8).isEmpty = '1') THEN
					addr_out <= store_buffer(8).address;
					opcode_out <= store_buffer(8).opcode;
					store_buffer(8).isEmpty <= '0';
				ELSIF(store_buffer(9).isEmpty = '1') THEN
					addr_out <= store_buffer(9).address;
					opcode_out <= store_buffer(9).opcode;
					store_buffer(9).isEmpty <= '0';
				ELSIF(store_buffer(10).isEmpty = '1') THEN
					addr_out <= store_buffer(10).address;
					opcode_out <= store_buffer(10).opcode;
					store_buffer(10).isEmpty <= '0';
				ELSIF(store_buffer(11).isEmpty = '1') THEN
					addr_out <= store_buffer(11).address;
					opcode_out <= store_buffer(11).opcode;
					store_buffer(11).isEmpty <= '0';
				ELSIF(store_buffer(12).isEmpty = '1') THEN
					addr_out <= store_buffer(12).address;
					opcode_out <= store_buffer(12).opcode;
					store_buffer(12).isEmpty <= '0';
				ELSIF(store_buffer(13).isEmpty = '1') THEN
					addr_out <= store_buffer(13).address;
					opcode_out <= store_buffer(13).opcode;
					store_buffer(13).isEmpty <= '0';
				ELSIF(store_buffer(14).isEmpty = '1') THEN
					addr_out <= store_buffer(14).address;
					opcode_out <= store_buffer(14).opcode;
					store_buffer(14).isEmpty <= '0';
				ELSIF(store_buffer(15).isEmpty = '1') THEN
					addr_out <= store_buffer(15).address;
					opcode_out <= store_buffer(15).opcode;
					store_buffer(15).isEmpty <= '0';
				ELSIF(store_buffer(16).isEmpty = '1') THEN
					addr_out <= store_buffer(16).address;
					opcode_out <= store_buffer(16).opcode;
					store_buffer(16).isEmpty <= '0';
				ELSIF(store_buffer(17).isEmpty = '1') THEN
					addr_out <= store_buffer(17).address;
					opcode_out <= store_buffer(17).opcode;
					store_buffer(17).isEmpty <= '0';
				ELSIF(store_buffer(18).isEmpty = '1') THEN
					addr_out <= store_buffer(18).address;
					opcode_out <= store_buffer(18).opcode;
					store_buffer(18).isEmpty <= '0';
				ELSIF(store_buffer(19).isEmpty = '1') THEN
					addr_out <= store_buffer(19).address;
					opcode_out <= store_buffer(19).opcode;
					store_buffer(19).isEmpty <= '0';
				ELSIF(store_buffer(20).isEmpty = '1') THEN
					addr_out <= store_buffer(20).address;
					opcode_out <= store_buffer(20).opcode;
					store_buffer(20).isEmpty <= '0';
				ELSIF(store_buffer(21).isEmpty = '1') THEN
					addr_out <= store_buffer(21).address;
					opcode_out <= store_buffer(21).opcode;
					store_buffer(21).isEmpty <= '0';
				ELSIF(store_buffer(22).isEmpty = '1') THEN
					addr_out <= store_buffer(22).address;
					opcode_out <= store_buffer(22).opcode;
					store_buffer(22).isEmpty <= '0';
				ELSIF(store_buffer(23).isEmpty = '1') THEN
					addr_out <= store_buffer(23).address;
					opcode_out <= store_buffer(23).opcode;
					store_buffer(23).isEmpty <= '0';
				ELSIF(store_buffer(24).isEmpty = '1') THEN
					addr_out <= store_buffer(24).address;
					opcode_out <= store_buffer(24).opcode;
					store_buffer(24).isEmpty <= '0';
				ELSIF(store_buffer(25).isEmpty = '1') THEN
					addr_out <= store_buffer(25).address;
					opcode_out <= store_buffer(25).opcode;
					store_buffer(25).isEmpty <= '0';
				ELSIF(store_buffer(26).isEmpty = '1') THEN
					addr_out <= store_buffer(26).address;
					opcode_out <= store_buffer(26).opcode;
					store_buffer(26).isEmpty <= '0';
				ELSIF(store_buffer(27).isEmpty = '1') THEN
					addr_out <= store_buffer(27).address;
					opcode_out <= store_buffer(27).opcode;
					store_buffer(27).isEmpty <= '0';
				ELSIF(store_buffer(28).isEmpty = '1') THEN
					addr_out <= store_buffer(28).address;
					opcode_out <= store_buffer(28).opcode;
					store_buffer(28).isEmpty <= '0';
				ELSIF(store_buffer(29).isEmpty = '1') THEN
					addr_out <= store_buffer(29).address;
					opcode_out <= store_buffer(29).opcode;
					store_buffer(29).isEmpty <= '0';
				ELSIF(store_buffer(30).isEmpty = '1') THEN
					addr_out <= store_buffer(30).address;
					opcode_out <= store_buffer(30).opcode;
					store_buffer(30).isEmpty <= '0';
				ELSIF(store_buffer(31).isEmpty = '1') THEN
					addr_out <= store_buffer(31).address;
					opcode_out <= store_buffer(31).opcode;
					store_buffer(31).isEmpty <= '0';
				END IF;
			ELSE
				store_in	<=	'0';
			END IF;
			---
			IF(store_buffer(0).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(1).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(1).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(2).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(3).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(4).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(5).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(6).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(7).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(8).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(9).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(10).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(11).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(12).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(13).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(14).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(15).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(16).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(17).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(18).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(19).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(20).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(21).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(22).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(23).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(24).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(25).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(26).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(27).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(28).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(29).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(30).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSIF(store_buffer(31).isEmpty = '1') THEN
				store_buff_empty_sig <= '0';
			ELSE
				store_buff_empty_sig <= '1';
			END IF;
			----
			IF(load_buffer(0).isEmpty = '0') THEN--load buffer full?
				load_buff_full <= '0';
			ELSIF(load_buffer(1).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(1).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(2).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(3).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(4).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(5).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(6).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(7).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(8).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(9).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(10).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(11).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(12).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(13).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(14).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(15).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(16).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(17).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(18).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(19).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(20).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(21).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(22).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(23).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(24).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(25).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(26).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(27).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(28).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(29).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(30).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSIF(load_buffer(31).isEmpty = '0') THEN
				load_buff_full <= '0';
			ELSE
				load_buff_full <= '1';
			END IF;
			----
			IF(store_buffer(0).isEmpty = '0') THEN--store buffer full?
				store_buff_full <= '0';
			ELSIF(store_buffer(1).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(1).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(2).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(3).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(4).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(5).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(6).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(7).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(8).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(9).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(10).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(11).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(12).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(13).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(14).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(15).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(16).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(17).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(18).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(19).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(20).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(21).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(22).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(23).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(24).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(25).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(26).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(27).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(28).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(29).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(30).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSIF(store_buffer(31).isEmpty = '0') THEN
				store_buff_full <= '0';
			ELSE
				store_buff_full <= '1';
			END IF;
			-----
			IF((MEM_busy = '0') AND (store_buff_empty_sig = '1')) THEN--pushing items into the mem unit
				load_in	<=	'1';
				IF(load_buffer(0).isEmpty = '1') THEN
					addr_out <= load_buffer(0).address;
					opcode_out <= load_buffer(0).opcode;
					load_buffer(0).isEmpty <= '0';
				ELSIF(load_buffer(1).isEmpty = '1') THEN
					addr_out <= load_buffer(1).address;
					opcode_out <= load_buffer(1).opcode;
					load_buffer(1).isEmpty <= '0';
				ELSIF(load_buffer(2).isEmpty = '1') THEN
					addr_out <= load_buffer(2).address;
					opcode_out <= load_buffer(2).opcode;
					load_buffer(2).isEmpty <= '0';
				ELSIF(load_buffer(3).isEmpty = '1') THEN
					addr_out <= load_buffer(3).address;
					opcode_out <= load_buffer(3).opcode;
					load_buffer(3).isEmpty <= '0';
				ELSIF(load_buffer(4).isEmpty = '1') THEN
					addr_out <= load_buffer(4).address;
					opcode_out <= load_buffer(4).opcode;
					load_buffer(4).isEmpty <= '0';
				ELSIF(load_buffer(5).isEmpty = '1') THEN
					addr_out <= load_buffer(5).address;
					opcode_out <= load_buffer(5).opcode;
					load_buffer(5).isEmpty <= '0';
				ELSIF(load_buffer(6).isEmpty = '1') THEN
					addr_out <= load_buffer(6).address;
					opcode_out <= load_buffer(6).opcode;
					load_buffer(6).isEmpty <= '0';
				ELSIF(load_buffer(7).isEmpty = '1') THEN
					addr_out <= load_buffer(7).address;
					opcode_out <= load_buffer(7).opcode;
					load_buffer(7).isEmpty <= '0';
				ELSIF(load_buffer(8).isEmpty = '1') THEN
					addr_out <= load_buffer(8).address;
					opcode_out <= load_buffer(8).opcode;
					load_buffer(8).isEmpty <= '0';
				ELSIF(load_buffer(9).isEmpty = '1') THEN
					addr_out <= load_buffer(9).address;
					opcode_out <= load_buffer(9).opcode;
					load_buffer(9).isEmpty <= '0';
				ELSIF(load_buffer(10).isEmpty = '1') THEN
					addr_out <= load_buffer(10).address;
					opcode_out <= load_buffer(10).opcode;
					load_buffer(10).isEmpty <= '0';
				ELSIF(load_buffer(11).isEmpty = '1') THEN
					addr_out <= load_buffer(11).address;
					opcode_out <= load_buffer(11).opcode;
					load_buffer(11).isEmpty <= '0';
				ELSIF(load_buffer(12).isEmpty = '1') THEN
					addr_out <= load_buffer(12).address;
					opcode_out <= load_buffer(12).opcode;
					load_buffer(12).isEmpty <= '0';
				ELSIF(load_buffer(13).isEmpty = '1') THEN
					addr_out <= load_buffer(13).address;
					opcode_out <= load_buffer(13).opcode;
					load_buffer(13).isEmpty <= '0';
				ELSIF(load_buffer(14).isEmpty = '1') THEN
					addr_out <= load_buffer(14).address;
					opcode_out <= load_buffer(14).opcode;
					load_buffer(14).isEmpty <= '0';
				ELSIF(load_buffer(15).isEmpty = '1') THEN
					addr_out <= load_buffer(15).address;
					opcode_out <= load_buffer(15).opcode;
					load_buffer(15).isEmpty <= '0';
				ELSIF(load_buffer(16).isEmpty = '1') THEN
					addr_out <= load_buffer(16).address;
					opcode_out <= load_buffer(16).opcode;
					load_buffer(16).isEmpty <= '0';
				ELSIF(load_buffer(17).isEmpty = '1') THEN
					addr_out <= load_buffer(17).address;
					opcode_out <= load_buffer(17).opcode;
					load_buffer(17).isEmpty <= '0';
				ELSIF(load_buffer(18).isEmpty = '1') THEN
					addr_out <= load_buffer(18).address;
					opcode_out <= load_buffer(18).opcode;
					load_buffer(18).isEmpty <= '0';
				ELSIF(load_buffer(19).isEmpty = '1') THEN
					addr_out <= load_buffer(19).address;
					opcode_out <= load_buffer(19).opcode;
					load_buffer(19).isEmpty <= '0';
				ELSIF(load_buffer(20).isEmpty = '1') THEN
					addr_out <= load_buffer(20).address;
					opcode_out <= load_buffer(20).opcode;
					load_buffer(20).isEmpty <= '0';
				ELSIF(load_buffer(21).isEmpty = '1') THEN
					addr_out <= load_buffer(21).address;
					opcode_out <= load_buffer(21).opcode;
					load_buffer(21).isEmpty <= '0';
				ELSIF(load_buffer(22).isEmpty = '1') THEN
					addr_out <= load_buffer(22).address;
					opcode_out <= load_buffer(22).opcode;
					load_buffer(22).isEmpty <= '0';
				ELSIF(load_buffer(23).isEmpty = '1') THEN
					addr_out <= load_buffer(23).address;
					opcode_out <= load_buffer(23).opcode;
					load_buffer(23).isEmpty <= '0';
				ELSIF(load_buffer(24).isEmpty = '1') THEN
					addr_out <= load_buffer(24).address;
					opcode_out <= load_buffer(24).opcode;
					load_buffer(24).isEmpty <= '0';
				ELSIF(load_buffer(25).isEmpty = '1') THEN
					addr_out <= load_buffer(25).address;
					opcode_out <= load_buffer(25).opcode;
					load_buffer(25).isEmpty <= '0';
				ELSIF(load_buffer(26).isEmpty = '1') THEN
					addr_out <= load_buffer(26).address;
					opcode_out <= load_buffer(26).opcode;
					load_buffer(26).isEmpty <= '0';
				ELSIF(load_buffer(27).isEmpty = '1') THEN
					addr_out <= load_buffer(27).address;
					opcode_out <= load_buffer(27).opcode;
					load_buffer(27).isEmpty <= '0';
				ELSIF(load_buffer(28).isEmpty = '1') THEN
					addr_out <= load_buffer(28).address;
					opcode_out <= load_buffer(28).opcode;
					load_buffer(28).isEmpty <= '0';
				ELSIF(load_buffer(29).isEmpty = '1') THEN
					addr_out <= load_buffer(29).address;
					opcode_out <= load_buffer(29).opcode;
					load_buffer(29).isEmpty <= '0';
				ELSIF(load_buffer(30).isEmpty = '1') THEN
					addr_out <= load_buffer(30).address;
					opcode_out <= load_buffer(30).opcode;
					load_buffer(30).isEmpty <= '0';
				ELSIF(load_buffer(31).isEmpty = '1') THEN
					addr_out <= load_buffer(31).address;
					opcode_out <= load_buffer(31).opcode;
					load_buffer(31).isEmpty <= '0';
				END IF;
			ELSE
				load_in	<=	'0';
			END IF;
			
			IF(MEM_busy = '1') THEN
				addr_out <= X"00000000";
				opcode_out <= "000000";
			END IF;
			
		END IF;
	END PROCESS;

END behavior;